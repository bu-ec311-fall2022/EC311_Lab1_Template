`timescale 1ns / 1ps

// EC-311 Lab-1 Part-1
  // The names of the variables are as described in the lab handout

module add_sub_4_bit #
(
  parameter WIDTH = 4
)
(
  // The inputs 
  input wire [WIDTH-1:0]        A_input,
  input wire [WIDTH-1:0]        B_input,
  input wire                    M_control_input,

  // The outputs
  output wire                   V_out,
  output wire                   C_out,
  output wire [WIDTH-1:0]       S_output

);



endmodule
